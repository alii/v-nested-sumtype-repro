module token

pub const keyword_map = {
	'fn': Kind.kw_function
}
