module flags

pub struct Flags {
pub:
	expose_debug_builtins bool
	io_enabled            bool
	std_lib_enabled       bool
}
