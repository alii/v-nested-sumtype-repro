module span

pub struct Span {
pub:
	start_line   int
	start_column int
	end_line     int
	end_column   int
}
